module full_adder_withoutC (input a, input b, input cin, output s);
    xor(s, a, b, cin);
endmodule
